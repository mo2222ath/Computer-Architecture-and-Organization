module Ex_34(
	Ta,
	Tb,
	Clk,
	La1,
	La0,
	Lb1,
	Lb0
);


input wire	Ta;
input wire	Tb;
input wire	Clk;
output wire	La1;
output wire	La0;
output wire	Lb1;
output wire	Lb0;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
reg	SYNTHESIZED_WIRE_11;
reg	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;

assign	La1 = SYNTHESIZED_WIRE_11;



assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_1;

assign	SYNTHESIZED_WIRE_3 =  ~SYNTHESIZED_WIRE_11;

assign	SYNTHESIZED_WIRE_4 =  ~SYNTHESIZED_WIRE_12;

assign	SYNTHESIZED_WIRE_5 =  ~Ta;

assign	SYNTHESIZED_WIRE_6 =  ~SYNTHESIZED_WIRE_11;

assign	Lb0 = SYNTHESIZED_WIRE_12 & SYNTHESIZED_WIRE_11;

assign	SYNTHESIZED_WIRE_7 =  ~SYNTHESIZED_WIRE_12;

assign	SYNTHESIZED_WIRE_8 =  ~Tb;

assign	La0 = SYNTHESIZED_WIRE_2 & SYNTHESIZED_WIRE_12;

assign	SYNTHESIZED_WIRE_1 = SYNTHESIZED_WIRE_3 & SYNTHESIZED_WIRE_4 & SYNTHESIZED_WIRE_5;

assign	SYNTHESIZED_WIRE_0 = SYNTHESIZED_WIRE_6 & SYNTHESIZED_WIRE_7 & SYNTHESIZED_WIRE_8;

assign	SYNTHESIZED_WIRE_10 = SYNTHESIZED_WIRE_11 ^ SYNTHESIZED_WIRE_12;

assign	SYNTHESIZED_WIRE_2 =  ~SYNTHESIZED_WIRE_11;

assign	Lb1 =  ~SYNTHESIZED_WIRE_11;


always@(posedge Clk)
begin
	begin
	SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_9;
	end
end

always@(posedge Clk)
begin
	begin
	SYNTHESIZED_WIRE_11 <= SYNTHESIZED_WIRE_10;
	end
end


endmodule
